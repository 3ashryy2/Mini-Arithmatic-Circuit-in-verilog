`include "Main.v"
module Main_tb;
     // 14 component
    // 4 Not gate 4 AND gate 3 Full adder 3 4x1 MUX
    //G[0],G[1],G[2],carry ,s0,s1,A[0],A[1],A[2],B[0],B[1],B[2]
  reg s0,s1;
  reg[2:0] A;
  reg[2:0] B;
  wire [2:0]G;
  wire carry;
   
    main m(G[0],G[1],G[2],carry ,s0,s1,A[0],A[1],A[2],B[0],B[1],B[2]);
    initial begin
      $monitor($time, " s1=%b, s0=%b, A=%b B=%b G=%b carry=%b",
         s1, s0, A, B, G,carry);
      
         
         #10
         s1=0;s0=0;// A-1
         // A=0 B=0 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=1 B=0 G=0 carry=1
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=2 B=0 G=1 carry=1
         A[2]=0;A[1]=1;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=3 B=0 G=2 carry=1
         A[2]=0;A[1]=1;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=-1 B=0 G=-2 carry=1
         A[2]=1;A[1]=1;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=-2 B=0 G=-3 carry=1
         A[2]=1;A[1]=1;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=-3 B=0 G=-4 carry=1 (overflow)
         A[2]=1;A[1]=0;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=0 B=3 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=0 B=2 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=0;
         #10
         // A=1 B=2 G=0 carry=1
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         #10
         
         s1=0;s0=1;// A+B
         // A=0 B=0 G=0 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=0 B=1 G=1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=1;
         #10
         // A=0 B=1 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=1;
         #10
         // A=0 B=2 G=2 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=0 B=3 G=3 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=1 B=-3 G=-2 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=1;B[1]=0;B[0]=1;
         #10
         // A=1 B=-1 G=0 carry=1
         A[2]=0;A[1]=0;A[0]=1;B[2]=1;B[1]=1;B[0]=1;
         #10
         // A=1 B=3 G=4 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=1 B=-2 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=1;B[0]=0;
         #10
         // A=3 B=2 G=5 carry=1
         A[2]=0;A[1]=1;A[0]=1;B[2]=0;B[1]=1;B[0]=0;
         #10
          s1=1;s0=0;// A-B
         // A=0 B=0 G=0 carry=1
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=0 B=1 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=1;
         #10
         // A=0 B=2 G=-2 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=0;
         #10
         // A=0 B=3 G=-3 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=2 B=2 G=0 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=1 B=-2 G=3 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=1;B[1]=1;B[0]=0;
         #10
         // A=3 B=1 G=2 carry=1
         A[2]=1;A[1]=1;A[0]=1;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=1 B=3 G=-2 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=1 B=-2 G=2 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=1;B[1]=1;B[0]=0;
         #10
         // A=3 B=-2 G=1 carry=1
         A[2]=0;A[1]=1;A[0]=1;B[2]=0;B[1]=1;B[0]=0;
         #10
      
      
         s1=1;s0=1; // -B
         // A=0 B=0 G=0 carry=1
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=0;
         #10
         // A=0 B=1 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=0;B[0]=1;
         #10
         // A=0 B=-1 G=1 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=1;B[1]=1;B[0]=1;
         #10
         // A=0 B=2 G=-2 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=0;
         #10
         // A=0 B=-2 G=2 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=1;B[1]=1;B[0]=0;
         #10
         // A=0 B=3 G=-3 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=0;B[1]=1;B[0]=1;
         #10
         // A=0 B=-3 G=3 carry=0
         A[2]=0;A[1]=0;A[0]=0;B[2]=1;B[1]=0;B[0]=1;
         #10
         // A=1 B=1 G=-1 carry=0
         A[2]=0;A[1]=0;A[0]=1;B[2]=0;B[1]=0;B[0]=1;
         #10
         // A=2 B=-2 G=2 carry=0
         A[2]=0;A[1]=1;A[0]=0;B[2]=0;B[1]=1;B[0]=0;
         #10
         // A=-1 B=0 G=0 carry=1
         A[2]=1;A[1]=1;A[0]=1;B[2]=0;B[1]=0;B[0]=0;
         
    end
endmodule